module top();
trior v;
endmodule
