module top();
tri0 v;
endmodule
