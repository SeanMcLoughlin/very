class test_cls;
    int prop_a;
    int prop_b;
endclass
