`include "header.sv"
module test; endmodule