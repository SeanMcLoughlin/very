// Header file for include test
`define HEADER_LOADED 1