module incomplete_test(input clk