module top();
time signed v;
endmodule
