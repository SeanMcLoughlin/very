module top();
tri v;
endmodule
