module test(input clk, output reg data); endmodule