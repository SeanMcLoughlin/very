module test_gt; assign c = a > b; endmodule
module test_lt; assign c = a < b; endmodule
module test_gte; assign c = a >= b; endmodule
module test_lte; assign c = a <= b; endmodule