module test(clk, reset); endmodule