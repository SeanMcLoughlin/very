/*
:name: asinh_function
:description: $asinh test
:tags: 20.8
:type: simulation elaboration parsing
*/
module top();
initial
$display("%f", $asinh(4));
endmodule
