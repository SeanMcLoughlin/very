module top ();
    bit [7:0] arr[10];
endmodule
