module test(clk, data);
    input wire clk;
    output reg data;
endmodule