/*
:name: sin_function
:description: $sin test
:tags: 20.8
:type: simulation elaboration parsing
*/
module top();
initial
$display("%f", $sin(4));
endmodule
