module top();
    class test_cls;
        local int a_loc = 21;
        protected int a_prot = 22;
        int a = 23;
    endclass
    test_cls obj;

    initial begin

    end
endmodule
