module top();
tri1 v;
endmodule
