module top();
supply0 v;
endmodule
