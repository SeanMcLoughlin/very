module top();
integer unsigned v;
endmodule
