module top();
shortint unsigned v;
endmodule
