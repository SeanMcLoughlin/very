module test(input [3:0] a, output [7:0] result);
    assign result = a * 2 + 1;
endmodule