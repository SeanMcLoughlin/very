module top(input a, input b);

wire #10 w;

assign w = a & b;

endmodule
