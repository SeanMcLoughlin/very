module top();
logic a, b, c;
always_comb begin
    c = a & b;
end
endmodule
