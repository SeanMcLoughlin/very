/*
:name: tan_function
:description: $tan test
:tags: 20.8
:type: simulation elaboration parsing
*/
module top();
initial
$display("%f", $tan(4));
endmodule
