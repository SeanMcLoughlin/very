module top();
wire [7:0] a = 8'b1101x001;
endmodule
