module top ();
    integer mem[2][];
endmodule
