module top();
time unsigned v;
endmodule
