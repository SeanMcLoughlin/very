class test_cls;
    local int x = 42;
endclass
