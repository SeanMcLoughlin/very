class child extends parent;
    int y;
endclass
