module empty; endmodule