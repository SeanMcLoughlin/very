module top();
bit signed v;
endmodule
