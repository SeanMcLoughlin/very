`define WIDTH 8
module test; assign result = `WIDTH; endmodule