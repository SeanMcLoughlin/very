module top();
    logic a, clk;
    global clocking @(posedge clk); endclocking
endmodule
