module top();
integer signed v;
endmodule
