module top();
wire a;
endmodule
