module test; assign = invalid; endmodule