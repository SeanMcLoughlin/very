/*
:name: cosh_function
:description: $cosh test
:tags: 20.8
:type: simulation elaboration parsing
*/
module top();
initial
$display("%f", $cosh(4));
endmodule
