module top();
supply1 v;
endmodule
