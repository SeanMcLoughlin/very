module top();
longint unsigned v;
endmodule
