/*
:name: cos_function
:description: $cos test
:tags: 20.8
:type: simulation elaboration parsing
*/
module top();
initial
$display("%f", $cos(4));
endmodule
