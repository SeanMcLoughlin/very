/*
:name: atan_function
:description: $atan test
:tags: 20.8
:type: simulation elaboration parsing
*/
module top();
initial
$display("%f", $atan(4));
endmodule
