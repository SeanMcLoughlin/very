module top();
logic clk;
endmodule
