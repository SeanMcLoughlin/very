/*
:name: tanh_function
:description: $tanh test
:tags: 20.8
:type: simulation elaboration parsing
*/
module top();
initial
$display("%f", $tanh(4));
endmodule
