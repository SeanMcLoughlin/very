module test; assign c = a == b; endmodule