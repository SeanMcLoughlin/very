module top();
wire [7:0] data;
endmodule
