module top();
int count;
endmodule
