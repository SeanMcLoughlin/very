module top();
union {
    bit [7:0] v1;
    bit [3:0] v2;
} un;
endmodule
