module top();
uwire v;
endmodule
