/*
:name: atanh_function
:description: $atanh test
:tags: 20.8
:type: simulation elaboration parsing
*/
module top();
initial
$display("%f", $atanh(4));
endmodule
