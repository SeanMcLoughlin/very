module top();
trireg v;
endmodule
