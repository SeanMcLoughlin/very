module test; assign result = a + b; endmodule