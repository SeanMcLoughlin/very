module test; assign result = (a + b) * c; endmodule