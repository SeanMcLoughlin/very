module top ();
    bit [7:0] arr[];
endmodule
