module top();
int unsigned v;
endmodule
