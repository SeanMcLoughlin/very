module test(input [3:0] a, output b);
    assign b = ~&a;
endmodule