/*
:name: acos_function
:description: $acos test
:tags: 20.8
:type: simulation elaboration parsing
*/
module top();
initial
$display("%f", $acos(4));
endmodule
