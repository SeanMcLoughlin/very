/*
:name: asin_function
:description: $asin test
:tags: 20.8
:type: simulation elaboration parsing
*/
module top();
initial
$display("%f", $asin(4));
endmodule
