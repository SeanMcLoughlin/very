module top();
wand v;
endmodule
