module test(input clk, output data); assign data = clk; endmodule