module test; assign result = 42 * 3; endmodule