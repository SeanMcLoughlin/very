module top();
logic a, b;
always @(a) begin
    b = a;
end
endmodule
