class test_cls;
    protected int x = 42;
endclass
