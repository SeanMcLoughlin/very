class test_cls;
    int x;
endclass
