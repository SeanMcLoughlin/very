module top();
wor v;
endmodule
