module top();
wire c;
final begin
    $display(c);
end
endmodule
