module test(input [3:0] a, output [7:0] b); endmodule