/*
:name: sinh_function
:description: $sinh test
:tags: 20.8
:type: simulation elaboration parsing
*/
module top();
initial
$display("%f", $sinh(4));
endmodule
