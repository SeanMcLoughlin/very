module first; endmodule
module second(input clk); endmodule