module top();
byte unsigned v;
endmodule
