/*
:name: acosh_function
:description: $acosh test
:tags: 20.8
:type: simulation elaboration parsing
*/
module top();
initial
$display("%f", $acosh(4));
endmodule
