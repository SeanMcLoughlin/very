module top();
triand v;
endmodule
