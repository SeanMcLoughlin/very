module test; assign c = a != 8'b1101z001; endmodule